module subKeys(
    input [63:0] key, 
    output [47:0] sk1, sk2, sk3, sk4, sk5, sk6, sk7, sk8, sk9, sk10, sk11, sk12, sk13, sk14, sk15, sk16 );


    // 56 bit permutated key based on PC-1   
									
									// 63 - PC-1 values 
									
	wire [55:0] keyplus =  {key[7], key[15], key[23], key[31], key[39], key[47], key[55], key[63], key[6], key[14], key[22], key[30], key[38], key[46], key[54], key[62], key[5], key[13], key[21], key[29], key[37], key[45], key[53], key[61], key[4], key[12], key[20], key[28],  key[1], key[9],  key[17], key[25], key[33], key[41], key[49], key[57], key[2], key[10], key[18], key[26], key[34], key[42], key[50], key[58], key[3], key[11], key[19], key[27], key[35], key[43], key[51], key[59], key[36], key[44], key[52], key[60]};								
									
	 wire [27:0] C1, C2, C3, C4, C5, C6, C7, C8, C9, C10, C11, C12, C13, C14, C15, C16;
	 wire [27:0] D1, D2, D3, D4, D5, D6, D7, D8, D9, D10, D11, D12, D13, D14, D15, D16;								


    // C0 and D0  (split into left and right)

    wire [27:0] C0 = {keyplus[55-:28]};
    wire [27:0] D0 = {keyplus[27:0]};

			// 27 - PC-2

			assign sk1 =  {C1[14], C1[11], C1[17], C1[4], C1[27], C1[23], C1[25], C1[0], C1[13], C1[22], C1[7], C1[18], C1[5], C1[9], C1[16], C1[24], C1[2], C1[20], C1[12], C1[21], C1[1], C1[8], C1[15], C1[26], D1[15], D1[4], D1[25], D1[19], D1[9], D1[1], D1[26], D1[16], D1[5], D1[11], D1[23], D1[8], D1[12], D1[7], D1[17], D1[0], D1[22], D1[3], D1[10], D1[14], D1[6], D1[20], D1[27], D1[24] };
			assign sk2 =  {C2[14], C2[11], C2[17], C2[4], C2[27], C2[23], C2[25], C2[0], C2[13], C2[22], C2[7], C2[18], C2[5], C2[9], C2[16], C2[24], C2[2], C2[20], C2[12], C2[21], C2[1], C2[8], C2[15], C2[26], D2[15], D2[4], D2[25], D2[19], D2[9], D2[1], D2[26], D2[16], D2[5], D2[11], D2[23], D2[8], D2[12], D2[7], D2[17], D2[0], D2[22], D2[3], D2[10], D2[14], D2[6], D2[20], D2[27], D2[24] };
			assign sk3 =  {C3[14], C3[11], C3[17], C3[4], C3[27], C3[23], C3[25], C3[0], C3[13], C3[22], C3[7], C3[18], C3[5], C3[9], C3[16], C3[24], C3[2], C3[20], C3[12], C3[21], C3[1], C3[8], C3[15], C3[26], D3[15], D3[4], D3[25], D3[19], D3[9], D3[1], D3[26], D3[16], D3[5], D3[11], D3[23], D3[8], D3[12], D3[7], D3[17], D3[0], D3[22], D3[3], D3[10], D3[14], D3[6], D3[20], D3[27], D3[24] };
			assign sk4 =  {C4[14], C4[11], C4[17], C4[4], C4[27], C4[23], C4[25], C4[0], C4[13], C4[22], C4[7], C4[18], C4[5], C4[9], C4[16], C4[24], C4[2], C4[20], C4[12], C4[21], C4[1], C4[8], C4[15], C4[26], D4[15], D4[4], D4[25], D4[19], D4[9], D4[1], D4[26], D4[16], D4[5], D4[11], D4[23], D4[8], D4[12], D4[7], D4[17], D4[0], D4[22], D4[3], D4[10], D4[14], D4[6], D4[20], D4[27], D4[24] };
			assign sk5 =  {C5[14], C5[11], C5[17], C5[4], C5[27], C5[23], C5[25], C5[0], C5[13], C5[22], C5[7], C5[18], C5[5], C5[9], C5[16], C5[24], C5[2], C5[20], C5[12], C5[21], C5[1], C5[8], C5[15], C5[26], D5[15], D5[4], D5[25], D5[19], D5[9], D5[1], D5[26], D5[16], D5[5], D5[11], D5[23], D5[8], D5[12], D5[7], D5[17], D5[0], D5[22], D5[3], D5[10], D5[14], D5[6], D5[20], D5[27], D5[24] };
			assign sk6 =  {C6[14], C6[11], C6[17], C6[4], C6[27], C6[23], C6[25], C6[0], C6[13], C6[22], C6[7], C6[18], C6[5], C6[9], C6[16], C6[24], C6[2], C6[20], C6[12], C6[21], C6[1], C6[8], C6[15], C6[26], D6[15], D6[4], D6[25], D6[19], D6[9], D6[1], D6[26], D6[16], D6[5], D6[11], D6[23], D6[8], D6[12], D6[7], D6[17], D6[0], D6[22], D6[3], D6[10], D6[14], D6[6], D6[20], D6[27], D6[24] };
			assign sk7 =  {C7[14], C7[11], C7[17], C7[4], C7[27], C7[23], C7[25], C7[0], C7[13], C7[22], C7[7], C7[18], C7[5], C7[9], C7[16], C7[24], C7[2], C7[20], C7[12], C7[21], C7[1], C7[8], C7[15], C7[26], D7[15], D7[4], D7[25], D7[19], D7[9], D7[1], D7[26], D7[16], D7[5], D7[11], D7[23], D7[8], D7[12], D7[7], D7[17], D7[0], D7[22], D7[3], D7[10], D7[14], D7[6], D7[20], D7[27], D7[24] };
			assign sk8 =  {C8[14], C8[11], C8[17], C8[4], C8[27], C8[23], C8[25], C8[0], C8[13], C8[22], C8[7], C8[18], C8[5], C8[9], C8[16], C8[24], C8[2], C8[20], C8[12], C8[21], C8[1], C8[8], C8[15], C8[26], D8[15], D8[4], D8[25], D8[19], D8[9], D8[1], D8[26], D8[16], D8[5], D8[11], D8[23], D8[8], D8[12], D8[7], D8[17], D8[0], D8[22], D8[3], D8[10], D8[14], D8[6], D8[20], D8[27], D8[24] };
			assign sk9 =  {C9[14], C9[11], C9[17], C9[4], C9[27], C9[23], C9[25], C9[0], C9[13], C9[22], C9[7], C9[18], C9[5], C9[9], C9[16], C9[24], C9[2], C9[20], C9[12], C9[21], C9[1], C9[8], C9[15], C9[26], D9[15], D9[4], D9[25], D9[19], D9[9], D9[1], D9[26], D9[16], D9[5], D9[11], D9[23], D9[8], D9[12], D9[7], D9[17], D9[0], D9[22], D9[3], D9[10], D9[14], D9[6], D9[20], D9[27], D9[24] };
			assign sk10 = {C10[14], C10[11], C10[17], C10[4], C10[27], C10[23], C10[25], C10[0], C10[13], C10[22], C10[7], C10[18], C10[5], C10[9], C10[16], C10[24], C10[2], C10[20], C10[12], C10[21], C10[1], C10[8], C10[15], C10[26], D10[15], D10[4], D10[25], D10[19], D10[9], D10[1], D10[26], D10[16], D10[5], D10[11], D10[23], D10[8], D10[12], D10[7], D10[17], D10[0], D10[22], D10[3], D10[10], D10[14], D10[6], D10[20], D10[27], D10[24] };
			assign sk11 = {C11[14], C11[11], C11[17], C11[4], C11[27], C11[23], C11[25], C11[0], C11[13], C11[22], C11[7], C11[18], C11[5], C11[9], C11[16], C11[24], C11[2], C11[20], C11[12], C11[21], C11[1], C11[8], C11[15], C11[26], D11[15], D11[4], D11[25], D11[19], D11[9], D11[1], D11[26], D11[16], D11[5], D11[11], D11[23], D11[8], D11[12], D11[7], D11[17], D11[0], D11[22], D11[3], D11[10], D11[14], D11[6], D11[20], D11[27], D11[24] };
			assign sk12 = {C12[14], C12[11], C12[17], C12[4], C12[27], C12[23], C12[25], C12[0], C12[13], C12[22], C12[7], C12[18], C12[5], C12[9], C12[16], C12[24], C12[2], C12[20], C12[12], C12[21], C12[1], C12[8], C12[15], C12[26], D12[15], D12[4], D12[25], D12[19], D12[9], D12[1], D12[26], D12[16], D12[5], D12[11], D12[23], D12[8], D12[12], D12[7], D12[17], D12[0], D12[22], D12[3], D12[10], D12[14], D12[6], D12[20], D12[27], D12[24] };
			assign sk13 = {C13[14], C13[11], C13[17], C13[4], C13[27], C13[23], C13[25], C13[0], C13[13], C13[22], C13[7], C13[18], C13[5], C13[9], C13[16], C13[24], C13[2], C13[20], C13[12], C13[21], C13[1], C13[8], C13[15], C13[26], D13[15], D13[4], D13[25], D13[19], D13[9], D13[1], D13[26], D13[16], D13[5], D13[11], D13[23], D13[8], D13[12], D13[7], D13[17], D13[0], D13[22], D13[3], D13[10], D13[14], D13[6], D13[20], D13[27], D13[24] };
			assign sk14 = {C14[14], C14[11], C14[17], C14[4], C14[27], C14[23], C14[25], C14[0], C14[13], C14[22], C14[7], C14[18], C14[5], C14[9], C14[16], C14[24], C14[2], C14[20], C14[12], C14[21], C14[1], C14[8], C14[15], C14[26], D14[15], D14[4], D14[25], D14[19], D14[9], D14[1], D14[26], D14[16], D14[5], D14[11], D14[23], D14[8], D14[12], D14[7], D14[17], D14[0], D14[22], D14[3], D14[10], D14[14], D14[6], D14[20], D14[27], D14[24] };
			assign sk15 = {C15[14], C15[11], C15[17], C15[4], C15[27], C15[23], C15[25], C15[0], C15[13], C15[22], C15[7], C15[18], C15[5], C15[9], C15[16], C15[24], C15[2], C15[20], C15[12], C15[21], C15[1], C15[8], C15[15], C15[26], D15[15], D15[4], D15[25], D15[19], D15[9], D15[1], D15[26], D15[16], D15[5], D15[11], D15[23], D15[8], D15[12], D15[7], D15[17], D15[0], D15[22], D15[3], D15[10], D15[14], D15[6], D15[20], D15[27], D15[24] };
			assign sk16 = {C16[14], C16[11], C16[17], C16[4], C16[27], C16[23], C16[25], C16[0], C16[13], C16[22], C16[7], C16[18], C16[5], C16[9], C16[16], C16[24], C16[2], C16[20], C16[12], C16[21], C16[1], C16[8], C16[15], C16[26], D16[15], D16[4], D16[25], D16[19], D16[9], D16[1], D16[26], D16[16], D16[5], D16[11], D16[23], D16[8], D16[12], D16[7], D16[17], D16[0], D16[22], D16[3], D16[10], D16[14], D16[6], D16[20], D16[27], D16[24]};
			

			s1 S_C0(C0, C1);
			s1 S_C1(C1, C2);
			s2 S_C2(C2, C3);
			s2 S_C3(C3, C4);
			s2 S_C4(C4, C5);
			s2 S_C5(C5, C6);
			s2 S_C6(C6, C7);
			s2 S_C7(C7, C8);
			s1 S_C8(C8, C9);
			s2 S_C9(C9, C10);
			s2 S_C10(C10, C11);
			s2 S_C11(C11, C12);
			s2 S_C12(C12, C13);
			s2 S_C13(C13, C14);
			s2 S_C14(C14, C15);
			s1 S_C15(C15, C16);
			
			s1 S_D0(D0, D1);
			s1 S_D1(D1, D2);
			s2 S_D2(D2, D3);
			s2 S_D3(D3, D4);
			s2 S_D4(D4, D5);
			s2 S_D5(D5, D6);
			s2 S_D6(D6, D7);
			s2 S_D7(D7, D8);
			s1 S_D8(D8, D9);
			s2 S_D9(D9, D10);
			s2 S_D10(D10, D11);
			s2 S_D11(D11, D12);
			s2 S_D12(D12, D13);
			s2 S_D13(D13, D14);
			s2 S_D14(D14, D15);
			s1 S_D15(D15, D16);
			

endmodule


module s1(
	input [27:0]sk,
	output reg [27:0] shift);
	always @ (*)
	begin
			shift = {sk[26:0], sk[27]};    // shift 1
	end
endmodule	
	
module s2(
	input [27:0]sk,
	output reg [27:0] shift);
	always @ (*)
	begin
			shift = {sk[25:0], sk[27:26]}; // shift 2
	end
endmodule		
